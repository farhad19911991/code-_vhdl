THIS IS VHDL
