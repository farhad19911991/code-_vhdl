THIS IS VHDL

library ieee;
