THIS IS VHDL

this sen.
  .
  .
  .
  .
  This is end of file.
