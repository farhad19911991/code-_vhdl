THIS IS VHDL
  .
  .
  .
  .
  This is end of file.
This is another mod. 
