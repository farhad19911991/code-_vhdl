THIS IS VHDL

this sen.
