THIS IS VHDL
  .
  .
  .
  .
  
