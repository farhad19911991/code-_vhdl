THIS IS VHDL
  .
  .
  .
  .
  This is end of file.
