THIS IS VHDL
  library ieee;

this sen.
  .
  .
  .
 .
  This is end of file.
This is another mod. 
# this is 32-bit ....
